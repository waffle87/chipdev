module model #() ();
endmodule
